VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_newmot
  CLASS BLOCK ;
  FOREIGN wrapped_newmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 296.000 25.350 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.420 300.000 1.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.620 300.000 79.820 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.100 300.000 87.300 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.260 300.000 95.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.740 300.000 102.940 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.900 300.000 111.100 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.380 300.000 118.580 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.540 300.000 126.740 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.020 300.000 134.220 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.900 300.000 9.100 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.820 300.000 158.020 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.300 300.000 165.500 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.460 300.000 173.660 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.940 300.000 181.140 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.100 300.000 189.300 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.580 300.000 196.780 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.740 300.000 204.940 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.220 300.000 212.420 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.380 300.000 220.580 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.860 300.000 228.060 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.020 300.000 236.220 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.500 300.000 243.700 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.660 300.000 251.860 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.300 300.000 267.500 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.940 300.000 283.140 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.700 300.000 32.900 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.180 300.000 40.380 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 300.000 48.540 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.820 300.000 56.020 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.980 300.000 64.180 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.460 300.000 71.660 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.180 300.000 6.380 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.380 300.000 84.580 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.540 300.000 92.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.020 300.000 100.220 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.180 300.000 108.380 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.660 300.000 115.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.820 300.000 124.020 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.300 300.000 131.500 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.460 300.000 139.660 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.940 300.000 147.140 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.100 300.000 155.300 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.340 300.000 14.540 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.580 300.000 162.780 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 300.000 170.940 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.220 300.000 178.420 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.380 300.000 186.580 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.020 300.000 202.220 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.500 300.000 209.700 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.660 300.000 217.860 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.140 300.000 225.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.300 300.000 233.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.820 300.000 22.020 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.940 300.000 249.140 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.580 300.000 264.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.060 300.000 272.260 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.220 300.000 280.420 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.700 300.000 287.900 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 294.860 300.000 296.060 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.980 300.000 30.180 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.460 300.000 37.660 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.620 300.000 45.820 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.100 300.000 53.300 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.260 300.000 61.460 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 67.740 300.000 68.940 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.460 300.000 3.660 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.660 300.000 81.860 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.820 300.000 90.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.300 300.000 97.500 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.460 300.000 105.660 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.940 300.000 113.140 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.100 300.000 121.300 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.580 300.000 128.780 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 135.740 300.000 136.940 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.220 300.000 144.420 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.380 300.000 152.580 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.860 300.000 160.060 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.020 300.000 168.220 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.500 300.000 175.700 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.140 300.000 191.340 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.300 300.000 199.500 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.780 300.000 206.980 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.940 300.000 215.140 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.420 300.000 222.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.580 300.000 230.780 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.100 300.000 19.300 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.220 300.000 246.420 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.700 300.000 253.900 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.860 300.000 262.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 300.000 269.540 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.500 300.000 277.700 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 283.980 300.000 285.180 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.140 300.000 293.340 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.260 300.000 27.460 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.740 300.000 34.940 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 41.900 300.000 43.100 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.380 300.000 50.580 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.540 300.000 58.740 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 296.000 294.450 300.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.580 300.000 298.780 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 296.000 298.130 300.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 0.000 2.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.770 0.000 54.330 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.370 0.000 58.930 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970 0.000 63.530 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.170 0.000 72.730 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 0.000 82.390 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 0.000 86.990 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 0.000 7.410 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 0.000 96.190 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 0.000 100.790 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.290 0.000 105.850 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 0.000 110.450 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.490 0.000 115.050 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 0.000 119.650 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 0.000 124.250 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 0.000 129.310 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 0.000 133.910 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 0.000 138.510 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.450 0.000 12.010 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 0.000 143.110 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.150 0.000 147.710 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 0.000 16.610 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 0.000 21.210 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 0.000 25.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 0.000 35.470 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.210 0.000 152.770 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 0.000 199.230 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 0.000 204.290 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.330 0.000 208.890 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 0.000 213.490 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.530 0.000 218.090 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 0.000 222.690 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 0.000 227.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.390 0.000 236.950 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 0.000 241.550 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.810 0.000 157.370 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.590 0.000 246.150 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 0.000 250.750 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 0.000 255.810 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.850 0.000 260.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 0.000 265.010 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.050 0.000 269.610 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 0.000 274.210 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 0.000 283.870 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 0.000 288.470 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 0.000 161.970 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.510 0.000 293.070 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 0.000 297.670 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.010 0.000 166.570 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 0.000 171.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.210 0.000 175.770 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 0.000 185.430 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 0.000 194.630 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.380 4.000 152.580 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.060 4.000 204.260 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.820 4.000 209.020 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.580 4.000 213.780 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.660 4.000 217.860 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.420 4.000 222.620 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.180 4.000 227.380 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.940 4.000 232.140 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.700 4.000 236.900 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.140 4.000 157.340 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.220 4.000 246.420 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.980 4.000 251.180 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.740 4.000 255.940 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.820 4.000 260.020 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.580 4.000 264.780 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.100 4.000 274.300 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.860 4.000 279.060 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.620 4.000 283.820 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.380 4.000 288.580 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.900 4.000 162.100 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.140 4.000 293.340 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.660 4.000 166.860 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.420 4.000 171.620 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.500 4.000 175.700 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.020 4.000 185.220 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.540 4.000 194.740 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 296.000 29.030 300.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 296.000 2.350 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 296.000 6.030 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 296.000 21.210 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 296.000 48.350 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 296.000 86.530 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 296.000 90.670 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.790 296.000 94.350 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 296.000 98.030 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.610 296.000 102.170 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.290 296.000 105.850 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 296.000 109.990 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 296.000 113.670 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 296.000 117.350 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 296.000 121.490 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 296.000 52.030 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.610 296.000 125.170 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.290 296.000 128.850 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 296.000 132.990 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 296.000 136.670 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 296.000 140.350 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.930 296.000 144.490 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.610 296.000 148.170 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 296.000 152.310 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 296.000 155.990 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.110 296.000 159.670 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 296.000 56.170 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 296.000 163.810 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.930 296.000 167.490 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.290 296.000 59.850 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970 296.000 63.530 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 296.000 67.670 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 296.000 71.350 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 296.000 75.030 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.610 296.000 79.170 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.290 296.000 82.850 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 296.000 13.850 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 296.000 171.170 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 296.000 209.810 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 296.000 213.490 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 296.000 217.630 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.750 296.000 221.310 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 296.000 224.990 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 296.000 229.130 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.250 296.000 232.810 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.930 296.000 236.490 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 296.000 240.630 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 296.000 244.310 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 296.000 175.310 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 296.000 247.990 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.570 296.000 252.130 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 296.000 255.810 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 296.000 259.950 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.070 296.000 263.630 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 296.000 267.310 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.890 296.000 271.450 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 296.000 275.130 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.250 296.000 278.810 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 296.000 282.950 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 296.000 178.990 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 296.000 286.630 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 296.000 182.670 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.250 296.000 186.810 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930 296.000 190.490 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.610 296.000 194.170 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 296.000 198.310 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 296.000 201.990 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.570 296.000 206.130 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.020 4.000 49.220 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.060 4.000 68.260 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.580 4.000 77.780 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.100 4.000 87.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.180 4.000 91.380 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.700 4.000 100.900 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.220 4.000 110.420 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.980 4.000 115.180 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.500 4.000 124.700 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.260 4.000 129.460 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.340 4.000 133.540 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.620 4.000 11.820 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.860 4.000 143.060 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.620 4.000 147.820 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.380 4.000 16.580 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.900 4.000 26.100 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.660 4.000 30.860 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.420 4.000 35.620 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.180 4.000 40.380 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 296.000 32.710 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.290 296.000 36.850 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.970 296.000 40.530 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 296.000 44.210 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 296.000 9.710 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.970 296.000 17.530 300.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 297.475 289.595 ;
      LAYER met1 ;
        RECT 1.910 10.640 298.010 289.980 ;
      LAYER met2 ;
        RECT 2.630 295.720 5.190 298.365 ;
        RECT 6.310 295.720 8.870 298.365 ;
        RECT 9.990 295.720 13.010 298.365 ;
        RECT 14.130 295.720 16.690 298.365 ;
        RECT 17.810 295.720 20.370 298.365 ;
        RECT 21.490 295.720 24.510 298.365 ;
        RECT 25.630 295.720 28.190 298.365 ;
        RECT 29.310 295.720 31.870 298.365 ;
        RECT 32.990 295.720 36.010 298.365 ;
        RECT 37.130 295.720 39.690 298.365 ;
        RECT 40.810 295.720 43.370 298.365 ;
        RECT 44.490 295.720 47.510 298.365 ;
        RECT 48.630 295.720 51.190 298.365 ;
        RECT 52.310 295.720 55.330 298.365 ;
        RECT 56.450 295.720 59.010 298.365 ;
        RECT 60.130 295.720 62.690 298.365 ;
        RECT 63.810 295.720 66.830 298.365 ;
        RECT 67.950 295.720 70.510 298.365 ;
        RECT 71.630 295.720 74.190 298.365 ;
        RECT 75.310 295.720 78.330 298.365 ;
        RECT 79.450 295.720 82.010 298.365 ;
        RECT 83.130 295.720 85.690 298.365 ;
        RECT 86.810 295.720 89.830 298.365 ;
        RECT 90.950 295.720 93.510 298.365 ;
        RECT 94.630 295.720 97.190 298.365 ;
        RECT 98.310 295.720 101.330 298.365 ;
        RECT 102.450 295.720 105.010 298.365 ;
        RECT 106.130 295.720 109.150 298.365 ;
        RECT 110.270 295.720 112.830 298.365 ;
        RECT 113.950 295.720 116.510 298.365 ;
        RECT 117.630 295.720 120.650 298.365 ;
        RECT 121.770 295.720 124.330 298.365 ;
        RECT 125.450 295.720 128.010 298.365 ;
        RECT 129.130 295.720 132.150 298.365 ;
        RECT 133.270 295.720 135.830 298.365 ;
        RECT 136.950 295.720 139.510 298.365 ;
        RECT 140.630 295.720 143.650 298.365 ;
        RECT 144.770 295.720 147.330 298.365 ;
        RECT 148.450 295.720 151.470 298.365 ;
        RECT 152.590 295.720 155.150 298.365 ;
        RECT 156.270 295.720 158.830 298.365 ;
        RECT 159.950 295.720 162.970 298.365 ;
        RECT 164.090 295.720 166.650 298.365 ;
        RECT 167.770 295.720 170.330 298.365 ;
        RECT 171.450 295.720 174.470 298.365 ;
        RECT 175.590 295.720 178.150 298.365 ;
        RECT 179.270 295.720 181.830 298.365 ;
        RECT 182.950 295.720 185.970 298.365 ;
        RECT 187.090 295.720 189.650 298.365 ;
        RECT 190.770 295.720 193.330 298.365 ;
        RECT 194.450 295.720 197.470 298.365 ;
        RECT 198.590 295.720 201.150 298.365 ;
        RECT 202.270 295.720 205.290 298.365 ;
        RECT 206.410 295.720 208.970 298.365 ;
        RECT 210.090 295.720 212.650 298.365 ;
        RECT 213.770 295.720 216.790 298.365 ;
        RECT 217.910 295.720 220.470 298.365 ;
        RECT 221.590 295.720 224.150 298.365 ;
        RECT 225.270 295.720 228.290 298.365 ;
        RECT 229.410 295.720 231.970 298.365 ;
        RECT 233.090 295.720 235.650 298.365 ;
        RECT 236.770 295.720 239.790 298.365 ;
        RECT 240.910 295.720 243.470 298.365 ;
        RECT 244.590 295.720 247.150 298.365 ;
        RECT 248.270 295.720 251.290 298.365 ;
        RECT 252.410 295.720 254.970 298.365 ;
        RECT 256.090 295.720 259.110 298.365 ;
        RECT 260.230 295.720 262.790 298.365 ;
        RECT 263.910 295.720 266.470 298.365 ;
        RECT 267.590 295.720 270.610 298.365 ;
        RECT 271.730 295.720 274.290 298.365 ;
        RECT 275.410 295.720 277.970 298.365 ;
        RECT 279.090 295.720 282.110 298.365 ;
        RECT 283.230 295.720 285.790 298.365 ;
        RECT 286.910 295.720 289.470 298.365 ;
        RECT 290.590 295.720 293.610 298.365 ;
        RECT 294.730 295.720 297.290 298.365 ;
        RECT 1.940 4.280 297.980 295.720 ;
        RECT 1.940 2.195 1.970 4.280 ;
        RECT 3.090 2.195 6.570 4.280 ;
        RECT 7.690 2.195 11.170 4.280 ;
        RECT 12.290 2.195 15.770 4.280 ;
        RECT 16.890 2.195 20.370 4.280 ;
        RECT 21.490 2.195 24.970 4.280 ;
        RECT 26.090 2.195 30.030 4.280 ;
        RECT 31.150 2.195 34.630 4.280 ;
        RECT 35.750 2.195 39.230 4.280 ;
        RECT 40.350 2.195 43.830 4.280 ;
        RECT 44.950 2.195 48.430 4.280 ;
        RECT 49.550 2.195 53.490 4.280 ;
        RECT 54.610 2.195 58.090 4.280 ;
        RECT 59.210 2.195 62.690 4.280 ;
        RECT 63.810 2.195 67.290 4.280 ;
        RECT 68.410 2.195 71.890 4.280 ;
        RECT 73.010 2.195 76.950 4.280 ;
        RECT 78.070 2.195 81.550 4.280 ;
        RECT 82.670 2.195 86.150 4.280 ;
        RECT 87.270 2.195 90.750 4.280 ;
        RECT 91.870 2.195 95.350 4.280 ;
        RECT 96.470 2.195 99.950 4.280 ;
        RECT 101.070 2.195 105.010 4.280 ;
        RECT 106.130 2.195 109.610 4.280 ;
        RECT 110.730 2.195 114.210 4.280 ;
        RECT 115.330 2.195 118.810 4.280 ;
        RECT 119.930 2.195 123.410 4.280 ;
        RECT 124.530 2.195 128.470 4.280 ;
        RECT 129.590 2.195 133.070 4.280 ;
        RECT 134.190 2.195 137.670 4.280 ;
        RECT 138.790 2.195 142.270 4.280 ;
        RECT 143.390 2.195 146.870 4.280 ;
        RECT 147.990 2.195 151.930 4.280 ;
        RECT 153.050 2.195 156.530 4.280 ;
        RECT 157.650 2.195 161.130 4.280 ;
        RECT 162.250 2.195 165.730 4.280 ;
        RECT 166.850 2.195 170.330 4.280 ;
        RECT 171.450 2.195 174.930 4.280 ;
        RECT 176.050 2.195 179.990 4.280 ;
        RECT 181.110 2.195 184.590 4.280 ;
        RECT 185.710 2.195 189.190 4.280 ;
        RECT 190.310 2.195 193.790 4.280 ;
        RECT 194.910 2.195 198.390 4.280 ;
        RECT 199.510 2.195 203.450 4.280 ;
        RECT 204.570 2.195 208.050 4.280 ;
        RECT 209.170 2.195 212.650 4.280 ;
        RECT 213.770 2.195 217.250 4.280 ;
        RECT 218.370 2.195 221.850 4.280 ;
        RECT 222.970 2.195 226.910 4.280 ;
        RECT 228.030 2.195 231.510 4.280 ;
        RECT 232.630 2.195 236.110 4.280 ;
        RECT 237.230 2.195 240.710 4.280 ;
        RECT 241.830 2.195 245.310 4.280 ;
        RECT 246.430 2.195 249.910 4.280 ;
        RECT 251.030 2.195 254.970 4.280 ;
        RECT 256.090 2.195 259.570 4.280 ;
        RECT 260.690 2.195 264.170 4.280 ;
        RECT 265.290 2.195 268.770 4.280 ;
        RECT 269.890 2.195 273.370 4.280 ;
        RECT 274.490 2.195 278.430 4.280 ;
        RECT 279.550 2.195 283.030 4.280 ;
        RECT 284.150 2.195 287.630 4.280 ;
        RECT 288.750 2.195 292.230 4.280 ;
        RECT 293.350 2.195 296.830 4.280 ;
        RECT 297.950 2.195 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.400 297.180 295.600 298.345 ;
        RECT 4.400 296.500 296.000 297.180 ;
        RECT 3.070 296.460 296.000 296.500 ;
        RECT 3.070 294.460 295.600 296.460 ;
        RECT 3.070 293.740 296.000 294.460 ;
        RECT 4.400 291.740 295.600 293.740 ;
        RECT 3.070 291.020 296.000 291.740 ;
        RECT 3.070 289.020 295.600 291.020 ;
        RECT 3.070 288.980 296.000 289.020 ;
        RECT 4.400 288.300 296.000 288.980 ;
        RECT 4.400 286.980 295.600 288.300 ;
        RECT 3.070 286.300 295.600 286.980 ;
        RECT 3.070 285.580 296.000 286.300 ;
        RECT 3.070 284.220 295.600 285.580 ;
        RECT 4.400 283.580 295.600 284.220 ;
        RECT 4.400 283.540 296.000 283.580 ;
        RECT 4.400 282.220 295.600 283.540 ;
        RECT 3.070 281.540 295.600 282.220 ;
        RECT 3.070 280.820 296.000 281.540 ;
        RECT 3.070 279.460 295.600 280.820 ;
        RECT 4.400 278.820 295.600 279.460 ;
        RECT 4.400 278.100 296.000 278.820 ;
        RECT 4.400 277.460 295.600 278.100 ;
        RECT 3.070 276.100 295.600 277.460 ;
        RECT 3.070 275.380 296.000 276.100 ;
        RECT 3.070 274.700 295.600 275.380 ;
        RECT 4.400 273.380 295.600 274.700 ;
        RECT 4.400 272.700 296.000 273.380 ;
        RECT 3.070 272.660 296.000 272.700 ;
        RECT 3.070 270.660 295.600 272.660 ;
        RECT 3.070 269.940 296.000 270.660 ;
        RECT 4.400 267.940 295.600 269.940 ;
        RECT 3.070 267.900 296.000 267.940 ;
        RECT 3.070 265.900 295.600 267.900 ;
        RECT 3.070 265.180 296.000 265.900 ;
        RECT 4.400 263.180 295.600 265.180 ;
        RECT 3.070 262.460 296.000 263.180 ;
        RECT 3.070 260.460 295.600 262.460 ;
        RECT 3.070 260.420 296.000 260.460 ;
        RECT 4.400 259.740 296.000 260.420 ;
        RECT 4.400 258.420 295.600 259.740 ;
        RECT 3.070 257.740 295.600 258.420 ;
        RECT 3.070 257.020 296.000 257.740 ;
        RECT 3.070 256.340 295.600 257.020 ;
        RECT 4.400 255.020 295.600 256.340 ;
        RECT 4.400 254.340 296.000 255.020 ;
        RECT 3.070 254.300 296.000 254.340 ;
        RECT 3.070 252.300 295.600 254.300 ;
        RECT 3.070 252.260 296.000 252.300 ;
        RECT 3.070 251.580 295.600 252.260 ;
        RECT 4.400 250.260 295.600 251.580 ;
        RECT 4.400 249.580 296.000 250.260 ;
        RECT 3.070 249.540 296.000 249.580 ;
        RECT 3.070 247.540 295.600 249.540 ;
        RECT 3.070 246.820 296.000 247.540 ;
        RECT 4.400 244.820 295.600 246.820 ;
        RECT 3.070 244.100 296.000 244.820 ;
        RECT 3.070 242.100 295.600 244.100 ;
        RECT 3.070 242.060 296.000 242.100 ;
        RECT 4.400 241.380 296.000 242.060 ;
        RECT 4.400 240.060 295.600 241.380 ;
        RECT 3.070 239.380 295.600 240.060 ;
        RECT 3.070 238.660 296.000 239.380 ;
        RECT 3.070 237.300 295.600 238.660 ;
        RECT 4.400 236.660 295.600 237.300 ;
        RECT 4.400 236.620 296.000 236.660 ;
        RECT 4.400 235.300 295.600 236.620 ;
        RECT 3.070 234.620 295.600 235.300 ;
        RECT 3.070 233.900 296.000 234.620 ;
        RECT 3.070 232.540 295.600 233.900 ;
        RECT 4.400 231.900 295.600 232.540 ;
        RECT 4.400 231.180 296.000 231.900 ;
        RECT 4.400 230.540 295.600 231.180 ;
        RECT 3.070 229.180 295.600 230.540 ;
        RECT 3.070 228.460 296.000 229.180 ;
        RECT 3.070 227.780 295.600 228.460 ;
        RECT 4.400 226.460 295.600 227.780 ;
        RECT 4.400 225.780 296.000 226.460 ;
        RECT 3.070 225.740 296.000 225.780 ;
        RECT 3.070 223.740 295.600 225.740 ;
        RECT 3.070 223.020 296.000 223.740 ;
        RECT 4.400 221.020 295.600 223.020 ;
        RECT 3.070 220.980 296.000 221.020 ;
        RECT 3.070 218.980 295.600 220.980 ;
        RECT 3.070 218.260 296.000 218.980 ;
        RECT 4.400 216.260 295.600 218.260 ;
        RECT 3.070 215.540 296.000 216.260 ;
        RECT 3.070 214.180 295.600 215.540 ;
        RECT 4.400 213.540 295.600 214.180 ;
        RECT 4.400 212.820 296.000 213.540 ;
        RECT 4.400 212.180 295.600 212.820 ;
        RECT 3.070 210.820 295.600 212.180 ;
        RECT 3.070 210.100 296.000 210.820 ;
        RECT 3.070 209.420 295.600 210.100 ;
        RECT 4.400 208.100 295.600 209.420 ;
        RECT 4.400 207.420 296.000 208.100 ;
        RECT 3.070 207.380 296.000 207.420 ;
        RECT 3.070 205.380 295.600 207.380 ;
        RECT 3.070 205.340 296.000 205.380 ;
        RECT 3.070 204.660 295.600 205.340 ;
        RECT 4.400 203.340 295.600 204.660 ;
        RECT 4.400 202.660 296.000 203.340 ;
        RECT 3.070 202.620 296.000 202.660 ;
        RECT 3.070 200.620 295.600 202.620 ;
        RECT 3.070 199.900 296.000 200.620 ;
        RECT 4.400 197.900 295.600 199.900 ;
        RECT 3.070 197.180 296.000 197.900 ;
        RECT 3.070 195.180 295.600 197.180 ;
        RECT 3.070 195.140 296.000 195.180 ;
        RECT 4.400 194.460 296.000 195.140 ;
        RECT 4.400 193.140 295.600 194.460 ;
        RECT 3.070 192.460 295.600 193.140 ;
        RECT 3.070 191.740 296.000 192.460 ;
        RECT 3.070 190.380 295.600 191.740 ;
        RECT 4.400 189.740 295.600 190.380 ;
        RECT 4.400 189.700 296.000 189.740 ;
        RECT 4.400 188.380 295.600 189.700 ;
        RECT 3.070 187.700 295.600 188.380 ;
        RECT 3.070 186.980 296.000 187.700 ;
        RECT 3.070 185.620 295.600 186.980 ;
        RECT 4.400 184.980 295.600 185.620 ;
        RECT 4.400 184.260 296.000 184.980 ;
        RECT 4.400 183.620 295.600 184.260 ;
        RECT 3.070 182.260 295.600 183.620 ;
        RECT 3.070 181.540 296.000 182.260 ;
        RECT 3.070 180.860 295.600 181.540 ;
        RECT 4.400 179.540 295.600 180.860 ;
        RECT 4.400 178.860 296.000 179.540 ;
        RECT 3.070 178.820 296.000 178.860 ;
        RECT 3.070 176.820 295.600 178.820 ;
        RECT 3.070 176.100 296.000 176.820 ;
        RECT 4.400 174.100 295.600 176.100 ;
        RECT 3.070 174.060 296.000 174.100 ;
        RECT 3.070 172.060 295.600 174.060 ;
        RECT 3.070 172.020 296.000 172.060 ;
        RECT 4.400 171.340 296.000 172.020 ;
        RECT 4.400 170.020 295.600 171.340 ;
        RECT 3.070 169.340 295.600 170.020 ;
        RECT 3.070 168.620 296.000 169.340 ;
        RECT 3.070 167.260 295.600 168.620 ;
        RECT 4.400 166.620 295.600 167.260 ;
        RECT 4.400 165.900 296.000 166.620 ;
        RECT 4.400 165.260 295.600 165.900 ;
        RECT 3.070 163.900 295.600 165.260 ;
        RECT 3.070 163.180 296.000 163.900 ;
        RECT 3.070 162.500 295.600 163.180 ;
        RECT 4.400 161.180 295.600 162.500 ;
        RECT 4.400 160.500 296.000 161.180 ;
        RECT 3.070 160.460 296.000 160.500 ;
        RECT 3.070 158.460 295.600 160.460 ;
        RECT 3.070 158.420 296.000 158.460 ;
        RECT 3.070 157.740 295.600 158.420 ;
        RECT 4.400 156.420 295.600 157.740 ;
        RECT 4.400 155.740 296.000 156.420 ;
        RECT 3.070 155.700 296.000 155.740 ;
        RECT 3.070 153.700 295.600 155.700 ;
        RECT 3.070 152.980 296.000 153.700 ;
        RECT 4.400 150.980 295.600 152.980 ;
        RECT 3.070 150.260 296.000 150.980 ;
        RECT 3.070 148.260 295.600 150.260 ;
        RECT 3.070 148.220 296.000 148.260 ;
        RECT 4.400 147.540 296.000 148.220 ;
        RECT 4.400 146.220 295.600 147.540 ;
        RECT 3.070 145.540 295.600 146.220 ;
        RECT 3.070 144.820 296.000 145.540 ;
        RECT 3.070 143.460 295.600 144.820 ;
        RECT 4.400 142.820 295.600 143.460 ;
        RECT 4.400 142.780 296.000 142.820 ;
        RECT 4.400 141.460 295.600 142.780 ;
        RECT 3.070 140.780 295.600 141.460 ;
        RECT 3.070 140.060 296.000 140.780 ;
        RECT 3.070 138.700 295.600 140.060 ;
        RECT 4.400 138.060 295.600 138.700 ;
        RECT 4.400 137.340 296.000 138.060 ;
        RECT 4.400 136.700 295.600 137.340 ;
        RECT 3.070 135.340 295.600 136.700 ;
        RECT 3.070 134.620 296.000 135.340 ;
        RECT 3.070 133.940 295.600 134.620 ;
        RECT 4.400 132.620 295.600 133.940 ;
        RECT 4.400 131.940 296.000 132.620 ;
        RECT 3.070 131.900 296.000 131.940 ;
        RECT 3.070 129.900 295.600 131.900 ;
        RECT 3.070 129.860 296.000 129.900 ;
        RECT 4.400 129.180 296.000 129.860 ;
        RECT 4.400 127.860 295.600 129.180 ;
        RECT 3.070 127.180 295.600 127.860 ;
        RECT 3.070 127.140 296.000 127.180 ;
        RECT 3.070 125.140 295.600 127.140 ;
        RECT 3.070 125.100 296.000 125.140 ;
        RECT 4.400 124.420 296.000 125.100 ;
        RECT 4.400 123.100 295.600 124.420 ;
        RECT 3.070 122.420 295.600 123.100 ;
        RECT 3.070 121.700 296.000 122.420 ;
        RECT 3.070 120.340 295.600 121.700 ;
        RECT 4.400 119.700 295.600 120.340 ;
        RECT 4.400 118.980 296.000 119.700 ;
        RECT 4.400 118.340 295.600 118.980 ;
        RECT 3.070 116.980 295.600 118.340 ;
        RECT 3.070 116.260 296.000 116.980 ;
        RECT 3.070 115.580 295.600 116.260 ;
        RECT 4.400 114.260 295.600 115.580 ;
        RECT 4.400 113.580 296.000 114.260 ;
        RECT 3.070 113.540 296.000 113.580 ;
        RECT 3.070 111.540 295.600 113.540 ;
        RECT 3.070 111.500 296.000 111.540 ;
        RECT 3.070 110.820 295.600 111.500 ;
        RECT 4.400 109.500 295.600 110.820 ;
        RECT 4.400 108.820 296.000 109.500 ;
        RECT 3.070 108.780 296.000 108.820 ;
        RECT 3.070 106.780 295.600 108.780 ;
        RECT 3.070 106.060 296.000 106.780 ;
        RECT 4.400 104.060 295.600 106.060 ;
        RECT 3.070 103.340 296.000 104.060 ;
        RECT 3.070 101.340 295.600 103.340 ;
        RECT 3.070 101.300 296.000 101.340 ;
        RECT 4.400 100.620 296.000 101.300 ;
        RECT 4.400 99.300 295.600 100.620 ;
        RECT 3.070 98.620 295.600 99.300 ;
        RECT 3.070 97.900 296.000 98.620 ;
        RECT 3.070 96.540 295.600 97.900 ;
        RECT 4.400 95.900 295.600 96.540 ;
        RECT 4.400 95.860 296.000 95.900 ;
        RECT 4.400 94.540 295.600 95.860 ;
        RECT 3.070 93.860 295.600 94.540 ;
        RECT 3.070 93.140 296.000 93.860 ;
        RECT 3.070 91.780 295.600 93.140 ;
        RECT 4.400 91.140 295.600 91.780 ;
        RECT 4.400 90.420 296.000 91.140 ;
        RECT 4.400 89.780 295.600 90.420 ;
        RECT 3.070 88.420 295.600 89.780 ;
        RECT 3.070 87.700 296.000 88.420 ;
        RECT 4.400 85.700 295.600 87.700 ;
        RECT 3.070 84.980 296.000 85.700 ;
        RECT 3.070 82.980 295.600 84.980 ;
        RECT 3.070 82.940 296.000 82.980 ;
        RECT 4.400 82.260 296.000 82.940 ;
        RECT 4.400 80.940 295.600 82.260 ;
        RECT 3.070 80.260 295.600 80.940 ;
        RECT 3.070 80.220 296.000 80.260 ;
        RECT 3.070 78.220 295.600 80.220 ;
        RECT 3.070 78.180 296.000 78.220 ;
        RECT 4.400 77.500 296.000 78.180 ;
        RECT 4.400 76.180 295.600 77.500 ;
        RECT 3.070 75.500 295.600 76.180 ;
        RECT 3.070 74.780 296.000 75.500 ;
        RECT 3.070 73.420 295.600 74.780 ;
        RECT 4.400 72.780 295.600 73.420 ;
        RECT 4.400 72.060 296.000 72.780 ;
        RECT 4.400 71.420 295.600 72.060 ;
        RECT 3.070 70.060 295.600 71.420 ;
        RECT 3.070 69.340 296.000 70.060 ;
        RECT 3.070 68.660 295.600 69.340 ;
        RECT 4.400 67.340 295.600 68.660 ;
        RECT 4.400 66.660 296.000 67.340 ;
        RECT 3.070 66.620 296.000 66.660 ;
        RECT 3.070 64.620 295.600 66.620 ;
        RECT 3.070 64.580 296.000 64.620 ;
        RECT 3.070 63.900 295.600 64.580 ;
        RECT 4.400 62.580 295.600 63.900 ;
        RECT 4.400 61.900 296.000 62.580 ;
        RECT 3.070 61.860 296.000 61.900 ;
        RECT 3.070 59.860 295.600 61.860 ;
        RECT 3.070 59.140 296.000 59.860 ;
        RECT 4.400 57.140 295.600 59.140 ;
        RECT 3.070 56.420 296.000 57.140 ;
        RECT 3.070 54.420 295.600 56.420 ;
        RECT 3.070 54.380 296.000 54.420 ;
        RECT 4.400 53.700 296.000 54.380 ;
        RECT 4.400 52.380 295.600 53.700 ;
        RECT 3.070 51.700 295.600 52.380 ;
        RECT 3.070 50.980 296.000 51.700 ;
        RECT 3.070 49.620 295.600 50.980 ;
        RECT 4.400 48.980 295.600 49.620 ;
        RECT 4.400 48.940 296.000 48.980 ;
        RECT 4.400 47.620 295.600 48.940 ;
        RECT 3.070 46.940 295.600 47.620 ;
        RECT 3.070 46.220 296.000 46.940 ;
        RECT 3.070 45.540 295.600 46.220 ;
        RECT 4.400 44.220 295.600 45.540 ;
        RECT 4.400 43.540 296.000 44.220 ;
        RECT 3.070 43.500 296.000 43.540 ;
        RECT 3.070 41.500 295.600 43.500 ;
        RECT 3.070 40.780 296.000 41.500 ;
        RECT 4.400 38.780 295.600 40.780 ;
        RECT 3.070 38.060 296.000 38.780 ;
        RECT 3.070 36.060 295.600 38.060 ;
        RECT 3.070 36.020 296.000 36.060 ;
        RECT 4.400 35.340 296.000 36.020 ;
        RECT 4.400 34.020 295.600 35.340 ;
        RECT 3.070 33.340 295.600 34.020 ;
        RECT 3.070 33.300 296.000 33.340 ;
        RECT 3.070 31.300 295.600 33.300 ;
        RECT 3.070 31.260 296.000 31.300 ;
        RECT 4.400 30.580 296.000 31.260 ;
        RECT 4.400 29.260 295.600 30.580 ;
        RECT 3.070 28.580 295.600 29.260 ;
        RECT 3.070 27.860 296.000 28.580 ;
        RECT 3.070 26.500 295.600 27.860 ;
        RECT 4.400 25.860 295.600 26.500 ;
        RECT 4.400 25.140 296.000 25.860 ;
        RECT 4.400 24.500 295.600 25.140 ;
        RECT 3.070 23.140 295.600 24.500 ;
        RECT 3.070 22.420 296.000 23.140 ;
        RECT 3.070 21.740 295.600 22.420 ;
        RECT 4.400 20.420 295.600 21.740 ;
        RECT 4.400 19.740 296.000 20.420 ;
        RECT 3.070 19.700 296.000 19.740 ;
        RECT 3.070 17.700 295.600 19.700 ;
        RECT 3.070 17.660 296.000 17.700 ;
        RECT 3.070 16.980 295.600 17.660 ;
        RECT 4.400 15.660 295.600 16.980 ;
        RECT 4.400 14.980 296.000 15.660 ;
        RECT 3.070 14.940 296.000 14.980 ;
        RECT 3.070 12.940 295.600 14.940 ;
        RECT 3.070 12.220 296.000 12.940 ;
        RECT 4.400 10.220 295.600 12.220 ;
        RECT 3.070 9.500 296.000 10.220 ;
        RECT 3.070 7.500 295.600 9.500 ;
        RECT 3.070 7.460 296.000 7.500 ;
        RECT 4.400 6.780 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.780 ;
        RECT 3.070 4.780 295.600 5.460 ;
        RECT 3.070 4.060 296.000 4.780 ;
        RECT 3.070 3.380 295.600 4.060 ;
        RECT 4.400 2.215 295.600 3.380 ;
      LAYER met4 ;
        RECT 84.935 42.335 97.440 240.545 ;
        RECT 99.840 42.335 174.240 240.545 ;
        RECT 176.640 42.335 251.040 240.545 ;
        RECT 253.440 42.335 278.465 240.545 ;
  END
END wrapped_newmot
END LIBRARY

